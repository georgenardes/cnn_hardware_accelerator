-- top entity